/*
###############################################################################
# Copyright (c) 2019, PulseRain Technology LLC 
#
# This program is distributed under a dual license: an open source license, 
# and a commercial license. 
# 
# The open source license under which this program is distributed is the 
# GNU Public License version 3 (GPLv3).
#
# And for those who want to use this program in ways that are incompatible
# with the GPLv3, PulseRain Technology LLC offers commercial license instead.
# Please contact PulseRain Technology LLC (www.pulserain.com) for more detail.
#
###############################################################################
*/

`ifndef SDRAM_CONTROLLER_SVH
`define SDRAM_CONTROLLER_SVH

parameter int 	SDRAM_ADDR_BITS = 22;
parameter int   SDRAM_CAS = 3;
parameter int   SDRAM_DATA_BITS = 32;
parameter int   SDRAM_BUS_BITS = 16;


`endif

